module range_check
    (input logic val, low, high, 
    output logic is_between);


endmodule: range_check

module offset_check
    (input logic val, low, delta,
    output logic is_between);

endmodule: offset_check